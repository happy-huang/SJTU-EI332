library verilog;
use verilog.vl_types.all;
entity decode2to4_vlg_vec_tst is
end decode2to4_vlg_vec_tst;
