module io_output( 
		addr,datain,write_io_enable,io_clk,out_port0,out_port1,out_port2,out_port3  );

	input  [31:0]  addr,datain;  
	input    write_io_enable,io_clk;  
	output  [31:0] out_port0,out_port1,out_port2, out_port3;    
	reg  [31:0] out_port0;  
	reg [31:0] out_port1;  
	reg [31:0] out_port2;
	reg [31:0] out_port3;
	
	always @ (posedge io_clk)  
	begin   
		if (write_io_enable == 1)    
			case (addr[7:2])     
				6'b101010: out_port0 = datain; // 80h
				6'b100001: out_port1 = datain; // 84h     
				6'b100010: out_port2 = datain; // 88h
			   6'b100011: out_port3 = datain; // 88h	
				//  more ports，可根据需要设计更多的输出端口 
			endcase
	end
endmodule
