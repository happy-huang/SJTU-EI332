library verilog;
use verilog.vl_types.all;
entity cpu_io_vlg_vec_tst is
end cpu_io_vlg_vec_tst;
