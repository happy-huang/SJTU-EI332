library verilog;
use verilog.vl_types.all;
entity counter18_vlg_tst is
end counter18_vlg_tst;
